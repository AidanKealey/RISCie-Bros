// Datapath

module Datapath ()

endmodule