// Datapath

module Datapath ()